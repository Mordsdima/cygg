module main

import toml
import os
import encoding.hex
import crypto.ed25519
import encoding.base64
import x.json2

fn miner() ! {
	// mut bc := Blockchain{}

	mut conf_file := 'config.toml'

	if 'CONFIG' in os.environ() {
		conf_file = os.environ()['CONFIG']
	}

	cnf := toml.parse_file(conf_file) or { panic(err) }

	mut private := ed25519.PrivateKey{}

	if cnf.value('wallet.privateseed') == toml.null {
		println('No wallet found')
		// private = hex.encode(bcrypt.generate_salt().bytes())
		_, private = ed25519.generate_key()!
		mut f := os.open_append(conf_file) or { panic(err) }
		f.write_string("\n\n# THIS PART IS AUTOGENERATED\n[wallet]\nprivateseed=\"${hex.encode(private.seed())}\"") or {
			panic(err)
		}
		f.close()
		println('New generated wallet! Keep your config in ABSOLUTE secret!')
		panic('Restart application.')
	} else {
		private = ed25519.new_key_from_seed(hex.decode(cnf.value('wallet.privateseed').string())!)
		// unsafe { C.memcpy(&private[0], &cnf.value('wallet.private').array()[0], 32) }
	}

	mut mepeer := MePeer{
		skey: private
		port: u16(cnf.value('peer.port').int())
	}

	mepeer.init()

	for s in cnf.value('bootstrap.peers').array() {
		mepeer.add_peer(s.string())!
	}
	if cnf.value('bootstrap.peers').array().len == 0 {
		panic('Cant work without bootstrap peers')
	}

	p := private.public_key()
	waddr := base64.encode(p)

	for {
		println('requesting..')
		// lets get the latest block in order to get prev
		l := mepeer.request_last_block()!
		d := mepeer.request_difficulty()!
		mut block := Block{
			data:         json2.encode(CoinbaseTransaction{
				@type: 'coinbase'
				rig:   'Official Miner; UNSTABLE'
				to:    waddr
			})
			prev:         l
			diff:         d
			generated_by: waddr
			version:      0
		}
		block.signit(private)!
		println('Mining block with difficulty ${d}')
		block.mine(d)
		println('Successfully mined!')
		mepeer.add_new_block(mut block, false, Peer{ pkey: p })!
		// mepeer.update() or { panic(err) }
	}
}
